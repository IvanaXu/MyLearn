library verilog;
use verilog.vl_types.all;
entity BIN_to_BCD_BIN_to_BCD_0 is
    port(
        un1_BIN_to_BCD_0: out    vl_logic_vector(3 downto 1);
        un1_BIN_to_BCD_0_1: out    vl_logic_vector(3 downto 0);
        Q_NS_0          : in     vl_logic_vector(7 downto 1)
    );
end BIN_to_BCD_BIN_to_BCD_0;
