library verilog;
use verilog.vl_types.all;
entity testbench is
    generic(
        DELY            : integer := 20
    );
end testbench;
