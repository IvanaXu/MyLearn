library verilog;
use verilog.vl_types.all;
entity textbench is
    generic(
        DELY            : integer := 20
    );
end textbench;
