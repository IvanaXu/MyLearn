library verilog;
use verilog.vl_types.all;
entity testbench161 is
    generic(
        clock_period    : integer := 20
    );
end testbench161;
