library verilog;
use verilog.vl_types.all;
entity paomadeng_paomadeng_1_2 is
    port(
        sel_0_c         : in     vl_logic_vector(1 downto 0);
        led_0_c         : out    vl_logic_vector(7 downto 0);
        rst_c           : in     vl_logic;
        rst_c_0         : in     vl_logic;
        clk_c           : in     vl_logic
    );
end paomadeng_paomadeng_1_2;
