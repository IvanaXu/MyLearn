library verilog;
use verilog.vl_types.all;
entity testbench is
    generic(
        Key_0           : string  := "Key_0";
        Key_1           : string  := "Key_1";
        Key_2           : string  := "Key_1";
        Key_3           : string  := "Key_3";
        Key_4           : string  := "Key_4";
        Key_5           : string  := "Key_5";
        Key_6           : string  := "Key_6";
        Key_7           : string  := "Key_7";
        Key_8           : string  := "Key_8";
        Key_9           : string  := "Key_9";
        Key_A           : string  := "Key_A";
        Key_B           : string  := "Key_B";
        Key_C           : string  := "Key_C";
        Key_D           : string  := "Key_D";
        Key_E           : string  := "Key_E";
        Key_F           : string  := "Key_F";
        None            : string  := "None"
    );
end testbench;
